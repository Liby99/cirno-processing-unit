module memory (
	input [7:0] mem_in,
	input [7:0] addr,
	input memory_w_en, memory_r_en,
	input clk,
	output logic[7:0] mem_out
);
	logic [255:0][7:0] core;

	always @(posedge clk) begin
		if (memory_r_en)
			mem_out <= core[addr];
		if (memory_w_en)
			core[addr] <= mem_in;
	end
	initial begin
mem[0] = 8'b01010101;
mem[1] = 8'b00000101;
mem[2] = 8'b10110101;
mem[3] = 8'b00000110;
mem[4] = 8'b11001010;
mem[5] = 8'b00000100;
mem[6] = 8'b11100111;
mem[7] = 8'b00000010;
mem[8] = 8'b10101000;
mem[9] = 8'b00000101;
mem[10] = 8'b00000000;
mem[11] = 8'b00000000;
mem[12] = 8'b00000000;
mem[13] = 8'b00000000;
mem[14] = 8'b00000000;
mem[15] = 8'b00000000;
mem[16] = 8'b00000000;
mem[17] = 8'b00000000;
mem[18] = 8'b00000000;
mem[19] = 8'b00000000;
mem[20] = 8'b00000000;
mem[21] = 8'b00000000;
mem[22] = 8'b00000000;
mem[23] = 8'b00000000;
mem[24] = 8'b00000000;
mem[25] = 8'b00000000;
mem[26] = 8'b00000000;
mem[27] = 8'b00000000;
mem[28] = 8'b00000000;
mem[29] = 8'b00000000;
mem[30] = 8'b00000000;
mem[31] = 8'b00000000;
mem[32] = 8'b00000000;
mem[33] = 8'b00000000;
mem[34] = 8'b00000000;
mem[35] = 8'b00000000;
mem[36] = 8'b00000000;
mem[37] = 8'b00000000;
mem[38] = 8'b00000000;
mem[39] = 8'b00000000;
mem[40] = 8'b00000000;
mem[41] = 8'b00000000;
mem[42] = 8'b00000000;
mem[43] = 8'b00000000;
mem[44] = 8'b00000000;
mem[45] = 8'b00000000;
mem[46] = 8'b00000000;
mem[47] = 8'b00000000;
mem[48] = 8'b00000000;
mem[49] = 8'b00000000;
mem[50] = 8'b00000000;
mem[51] = 8'b00000000;
mem[52] = 8'b00000000;
mem[53] = 8'b00000000;
mem[54] = 8'b00000000;
mem[55] = 8'b00000000;
mem[56] = 8'b00000000;
mem[57] = 8'b00000000;
mem[58] = 8'b00000000;
mem[59] = 8'b00000000;
mem[60] = 8'b00000000;
mem[61] = 8'b00000000;
mem[62] = 8'b00000000;
mem[63] = 8'b00000000;
mem[64] = 8'b00000000;
mem[65] = 8'b00000000;
mem[66] = 8'b00000000;
mem[67] = 8'b00000000;
mem[68] = 8'b00000000;
mem[69] = 8'b00000000;
mem[70] = 8'b00000000;
mem[71] = 8'b00000000;
mem[72] = 8'b00000000;
mem[73] = 8'b00000000;
mem[74] = 8'b00000000;
mem[75] = 8'b00000000;
mem[76] = 8'b00000000;
mem[77] = 8'b00000000;
mem[78] = 8'b00000000;
mem[79] = 8'b00000000;
mem[80] = 8'b00000000;
mem[81] = 8'b00000000;
mem[82] = 8'b00000000;
mem[83] = 8'b00000000;
mem[84] = 8'b00000000;
mem[85] = 8'b00000000;
mem[86] = 8'b00000000;
mem[87] = 8'b00000000;
mem[88] = 8'b00000000;
mem[89] = 8'b00000000;
mem[90] = 8'b00000000;
mem[91] = 8'b00000000;
mem[92] = 8'b00000000;
mem[93] = 8'b00000000;
mem[94] = 8'b00000000;
mem[95] = 8'b00000000;
mem[96] = 8'b00000000;
mem[97] = 8'b00000000;
mem[98] = 8'b00000000;
mem[99] = 8'b00000000;
mem[100] = 8'b00000000;
mem[101] = 8'b00000000;
mem[102] = 8'b00000000;
mem[103] = 8'b00000000;
mem[104] = 8'b00000000;
mem[105] = 8'b00000000;
mem[106] = 8'b00000000;
mem[107] = 8'b00000000;
mem[108] = 8'b00000000;
mem[109] = 8'b00000000;
mem[110] = 8'b00000000;
mem[111] = 8'b00000000;
mem[112] = 8'b00000000;
mem[113] = 8'b00000000;
mem[114] = 8'b00000000;
mem[115] = 8'b00000000;
mem[116] = 8'b00000000;
mem[117] = 8'b00000000;
mem[118] = 8'b00000000;
mem[119] = 8'b00000000;
mem[120] = 8'b00000000;
mem[121] = 8'b00000000;
mem[122] = 8'b00000000;
mem[123] = 8'b00000000;
mem[124] = 8'b00000000;
mem[125] = 8'b00000000;
mem[126] = 8'b00000000;
mem[127] = 8'b00000000;
mem[128] = 8'b00000000;
mem[129] = 8'b00000000;
mem[130] = 8'b00000000;
mem[131] = 8'b00000000;
mem[132] = 8'b00000000;
mem[133] = 8'b00000000;
mem[134] = 8'b00000000;
mem[135] = 8'b00000000;
mem[136] = 8'b00000000;
mem[137] = 8'b00000000;
mem[138] = 8'b00000000;
mem[139] = 8'b00000000;
mem[140] = 8'b00000000;
mem[141] = 8'b00000000;
mem[142] = 8'b00000000;
mem[143] = 8'b00000000;
mem[144] = 8'b00000000;
mem[145] = 8'b00000000;
mem[146] = 8'b00000000;
mem[147] = 8'b00000000;
mem[148] = 8'b00000000;
mem[149] = 8'b00000000;
mem[150] = 8'b00000000;
mem[151] = 8'b00000000;
mem[152] = 8'b00000000;
mem[153] = 8'b00000000;
mem[154] = 8'b00000000;
mem[155] = 8'b00000000;
mem[156] = 8'b00000000;
mem[157] = 8'b00000000;
mem[158] = 8'b00000000;
mem[159] = 8'b00000000;
mem[160] = 8'b00000000;
mem[161] = 8'b00000000;
mem[162] = 8'b00000000;
mem[163] = 8'b00000000;
mem[164] = 8'b00000000;
mem[165] = 8'b00000000;
mem[166] = 8'b00000000;
mem[167] = 8'b00000000;
mem[168] = 8'b00000000;
mem[169] = 8'b00000000;
mem[170] = 8'b00000000;
mem[171] = 8'b00000000;
mem[172] = 8'b00000000;
mem[173] = 8'b00000000;
mem[174] = 8'b00000000;
mem[175] = 8'b00000000;
mem[176] = 8'b00000000;
mem[177] = 8'b00000000;
mem[178] = 8'b00000000;
mem[179] = 8'b00000000;
mem[180] = 8'b00000000;
mem[181] = 8'b00000000;
mem[182] = 8'b00000000;
mem[183] = 8'b00000000;
mem[184] = 8'b00000000;
mem[185] = 8'b00000000;
mem[186] = 8'b00000000;
mem[187] = 8'b00000000;
mem[188] = 8'b00000000;
mem[189] = 8'b00000000;
mem[190] = 8'b00000000;
mem[191] = 8'b00000000;
mem[192] = 8'b00000000;
mem[193] = 8'b00000000;
mem[194] = 8'b00000000;
mem[195] = 8'b00000000;
mem[196] = 8'b00000000;
mem[197] = 8'b00000000;
mem[198] = 8'b00000000;
mem[199] = 8'b00000000;
mem[200] = 8'b00000000;
mem[201] = 8'b00000000;
mem[202] = 8'b00000000;
mem[203] = 8'b00000000;
mem[204] = 8'b00000000;
mem[205] = 8'b00000000;
mem[206] = 8'b00000000;
mem[207] = 8'b00000000;
mem[208] = 8'b00000000;
mem[209] = 8'b00000000;
mem[210] = 8'b00000000;
mem[211] = 8'b00000000;
mem[212] = 8'b00000000;
mem[213] = 8'b00000000;
mem[214] = 8'b00000000;
mem[215] = 8'b00000000;
mem[216] = 8'b00000000;
mem[217] = 8'b00000000;
mem[218] = 8'b00000000;
mem[219] = 8'b00000000;
mem[220] = 8'b00000000;
mem[221] = 8'b00000000;
mem[222] = 8'b00000000;
mem[223] = 8'b00000000;
mem[224] = 8'b00000000;
mem[225] = 8'b00000000;
mem[226] = 8'b00000000;
mem[227] = 8'b00000000;
mem[228] = 8'b00000000;
mem[229] = 8'b00000000;
mem[230] = 8'b00000000;
mem[231] = 8'b00000000;
mem[232] = 8'b00000000;
mem[233] = 8'b00000000;
mem[234] = 8'b00000000;
mem[235] = 8'b00000000;
mem[236] = 8'b00000000;
mem[237] = 8'b00000000;
mem[238] = 8'b00000000;
mem[239] = 8'b00000000;
mem[240] = 8'b00000000;
mem[241] = 8'b00000000;
mem[242] = 8'b00000000;
mem[243] = 8'b00000000;
mem[244] = 8'b00000000;
mem[245] = 8'b00000000;
mem[246] = 8'b00000000;
mem[247] = 8'b00000000;
mem[248] = 8'b00000000;
mem[249] = 8'b00000000;
mem[250] = 8'b00000000;
mem[251] = 8'b00000000;
mem[252] = 8'b00000000;
mem[253] = 8'b00000000;
mem[254] = 8'b00000000;
mem[255] = 8'b00000000;

	end
endmodule
